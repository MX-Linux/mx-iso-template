   1)  Standard
   2)  persist_all     Snabb. Sparar root och home (använder RAM, spara vid avstängning)
   3)  persist_root    Snabb. Sparar enbart root (använder RAM, sparar vid avstängning)
   4)  persist_static  Långsam. Sparar root och home (ingen RAM-användning, sparar alltid)
   5)  persist_home    Bara home-persistens
   6)  frugal_persist  Frugal med både root och home-persistens
   7)  frugal_root     Frugal med enbart root persistens
   8)  frugal_static   Frugal med home och statisk root-persistens
   9)  frugal_home     Frugal med endast home-persistens
  10)  frugal_only     Bara Frugal, ingen persistens
