   1)  Standard
   2)  checkmd5        Kontrollera live-mediums integritet
   3)  checkfs         Kontrollera LiveUSB och persistens ext2/3/4 filsystem
   4)  toram           Kopiera det komprimerade filsystemet till RAM
   5)  from=usb        Slutför start från en LiveUSB
   6)  from=hd         Slutför start från en hårddisk
   7)  nousb2          Koppla från alla usb-2 enheter vid start
   8)  hwclock=ask     Få hjälp av systemet att avgöra klockans inställning
   9)  hwclock=utc     Hårdvaru-klockan använder UTC (Endast Linuxsystem)
  10)  hwclock=local   Hårdvaru-klocka använder lokal tid (Windows system)
  11)  password        Ändra lösenord före start
  12)  nostore         Stäng av LiveUSB-lagringsfunktionen (Endast LiveUSB)
  13)  dostore         Använd LiveUSB-lagringsfunktionen (Endast LiveUSB)
  14)  savestate       Spara en del filer vid omstarter (Endast LiveUSB)
  15)  nosavestate     Spara inte filer vid omstarter (Endast LiveUSB)
